//Definicion del modulo y su entradas y salidas
//Dentro del parentesis se definen las entradas y salidas 


module _and(input a, input b, output c);
//2.Definen cables o componentes internos 
//NA
//3. Asignaciones, instancias, conexiones

assign  c= a & b;
endmodule